library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY xUDP is 
	port(
		);
end xUDP;

ARCHITECTURE Structural of xUDP is

BEGIN

END Structural;